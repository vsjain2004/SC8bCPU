module IMEM_PRGM(A, B, C, D, E, F, G, H, I, J, K, L, M, N, O, P);
	output [15:0] A, B, C, D, E, F, G, H, I, J, K, L, M, N, O, P;
// add1
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001000000000100;
//	assign C = 16'b0011000000001011;
//	assign D = 16'b1111000000000000;
//	assign E = 16'b0000000000000000;
//	assign F = 16'b0000000000000000;
//	assign G = 16'b0000000000000000;
//	assign H = 16'b0000000000000000;
//	assign I = 16'b0000000000000000;
//	assign J = 16'b0000000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;
	
// add2	
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001010100000000;
//	assign C = 16'b0011010100000010;
//	assign D = 16'b1111000000000000;
//	assign E = 16'b0000000000000000;
//	assign F = 16'b0000000000000000;
//	assign G = 16'b0000000000000000;
//	assign H = 16'b0000000000000000;
//	assign I = 16'b0000000000000000;
//	assign J = 16'b0000000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;
	
//	add3
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001001100000100;
//	assign C = 16'b0101001100000000;
//	assign D = 16'b1111000000000000;
//	assign E = 16'b0000000000000000;
//	assign F = 16'b0000000000000000;
//	assign G = 16'b0000000000000000;
//	assign H = 16'b0000000000000000;
//	assign I = 16'b0000000000000000;
//	assign J = 16'b0000000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;

// add4
	assign A = 16'b0000000000000000;
	assign B = 16'b0001010000000000;
	assign C = 16'b0011100000000010;
	assign D = 16'b0000110000000000;
	assign E = 16'b0000000000000000;
	assign F = 16'b0000000000000000;
	assign G = 16'b0000000000000000;
	assign H = 16'b0000000000000000;
	assign I = 16'b0000000000000000;
	assign J = 16'b0000000000000000;
	assign K = 16'b0000000000000000;
	assign L = 16'b0000000000000000;
	assign M = 16'b0000000000000000;
	assign N = 16'b0000000000000000;
	assign O = 16'b0000000000000000;
	assign P = 16'b0000000000000000;

// add5	
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001010000000000;
//	assign C = 16'b0001001100000100;
//	assign D = 16'b0011110000000010;
//	assign E = 16'b1111000000000000;
//	assign F = 16'b0000000000000000;
//	assign G = 16'b0000000000000000;
//	assign H = 16'b0000000000000000;
//	assign I = 16'b0000000000000000;
//	assign J = 16'b0000000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;

// sub1
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001001000000100;
//	assign C = 16'b0100001000000010;
//	assign D = 16'b1111000000000000;
//	assign E = 16'b0000000000000000;
//	assign F = 16'b0000000000000000;
//	assign G = 16'b0000000000000000;
//	assign H = 16'b0000000000000000;
//	assign I = 16'b0000000000000000;
//	assign J = 16'b0000000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;
	
// sub2
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001010000000001;
//	assign C = 16'b0100010000000100;
//	assign D = 16'b1111000000000000;
//	assign E = 16'b0000000000000000;
//	assign F = 16'b0000000000000000;
//	assign G = 16'b0000000000000000;
//	assign H = 16'b0000000000000000;
//	assign I = 16'b0000000000000000;
//	assign J = 16'b0000000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;
	
// mul
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001000000000000;
//	assign C = 16'b0110001100000000;
//	assign D = 16'b0001010000000000;
//	assign E = 16'b0011010000000000;
//	assign F = 16'b0101001100000000;
//	assign G = 16'b1001011100000011;
//	assign H = 16'b1011000000000100;
//	assign I = 16'b0010010000000000;
//	assign J = 16'b1111000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;
	
// int div
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001001111111111;
//	assign C = 16'b0001010000000000;
//	assign D = 16'b0101001100000000;
//	assign E = 16'b0100010000000001;
//	assign F = 16'b0110000100000000;
//	assign G = 16'b1100000110000000;
//	assign H = 16'b1001000110000000;
//	assign I = 16'b1011000000000011;
//	assign J = 16'b1111000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;
	
// array traversal	
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001001100000000;
//	assign C = 16'b0001110000000000;
//	assign D = 16'b0101001100000000;
//	assign E = 16'b1001001100001000;
//	assign F = 16'b1011000000000010;
//	assign G = 16'b1111000000000000;
//	assign H = 16'b0000000000000000;
//	assign I = 16'b0000000000000000;
//	assign J = 16'b0000000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;
	
// cs1
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001010000000000;
//	assign C = 16'b1100000000000000;
//	assign D = 16'b0010010000000000;
//	assign E = 16'b0001001100000001;
//	assign F = 16'b0111000000000000;
//	assign G = 16'b0010110000000000;
//	assign H = 16'b0001010000000000;
//	assign I = 16'b1101000000000001;
//	assign J = 16'b0010010000000000;
//	assign K = 16'b1101000001111111;
//	assign L = 16'b0010010000000000;
//	assign M = 16'b1001000001111111;
//	assign N = 16'b1011000000001111;
//	assign O = 16'b1110000010000000;
//	assign P = 16'b1111000000000000;
	
// cs2
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001001100000000;
//	assign C = 16'b0001010000000000;
//	assign D = 16'b1100010000000001;
//	assign E = 16'b1001000000000000;
//	assign F = 16'b1011100000000111;
//	assign G = 16'b0101001100000000;
//	assign H = 16'b0001010000000001;
//	assign I = 16'b1001000000001000;
//	assign J = 16'b1011100000001101;
//	assign K = 16'b0011010000000001;
//	assign L = 16'b0010010000000001;
//	assign M = 16'b1010000000000010;
//	assign N = 16'b1111000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;

// countup
//	assign A = 16'b0000000000000000;
//	assign B = 16'b0001000011110101;
//	assign C = 16'b0101000000000000;
//	assign D = 16'b1000000000000000;
//	assign E = 16'b1001000000001010;
//	assign F = 16'b1011000000000010;
//	assign G = 16'b1111000000000000;
//	assign H = 16'b0000000000000000;
//	assign I = 16'b0000000000000000;
//	assign J = 16'b0000000000000000;
//	assign K = 16'b0000000000000000;
//	assign L = 16'b0000000000000000;
//	assign M = 16'b0000000000000000;
//	assign N = 16'b0000000000000000;
//	assign O = 16'b0000000000000000;
//	assign P = 16'b0000000000000000;
endmodule