module OR_5_bit(In1, In2, In3, In4, In5, Out);
	input In1, In2, In3, In4, In5;
	output Out;
	
	or(Out, In1, In2, In3, In4, In5);
	
endmodule