module busmux_4_to_1(In1, In2, In3, In4, s1, s0, Out);
	input [7:0] In1;
	input [7:0] In2;
	input [7:0] In3;
	input [7:0] In4;
	input s1, s0;
	output reg [7:0] Out;
	
	always@*
	begin
		case({s1, s0})
			2'b00: Out=In1;
			2'b01: Out=In2;
			2'b10: Out=In3;
			2'b11: Out=In4;
		endcase
	end
	
endmodule