module decoder5to32(S, O);
	input [4:0] S;
	output reg [31:0] O;
	
	always @(S)
	begin
		O = 32'b0;
		case({S})
			5'b00000: O[0]=1'b1;
			5'b00001: O[1]=1'b1;
			5'b00010: O[2]=1'b1;
			5'b00011: O[3]=1'b1;
			5'b00100: O[4]=1'b1;
			5'b00101: O[5]=1'b1;
			5'b00110: O[6]=1'b1;
			5'b00111: O[7]=1'b1;
			5'b01000: O[8]=1'b1;
			5'b01001: O[9]=1'b1;
			5'b01010: O[10]=1'b1;
			5'b01011: O[11]=1'b1;
			5'b01100: O[12]=1'b1;
			5'b01101: O[13]=1'b1;
			5'b01110: O[14]=1'b1;
			5'b01111: O[15]=1'b1;
			5'b10000: O[16]=1'b1;
			5'b10001: O[17]=1'b1;
			5'b10010: O[18]=1'b1;
			5'b10011: O[19]=1'b1;
			5'b10100: O[20]=1'b1;
			5'b10101: O[21]=1'b1;
			5'b10110: O[22]=1'b1;
			5'b10111: O[23]=1'b1;
			5'b11000: O[24]=1'b1;
			5'b11001: O[25]=1'b1;
			5'b11010: O[26]=1'b1;
			5'b11011: O[27]=1'b1;
			5'b11100: O[28]=1'b1;
			5'b11101: O[29]=1'b1;
			5'b11110: O[30]=1'b1;
			5'b11111: O[31]=1'b1;
		endcase
	end
endmodule