module decoder4to16(S, O);
	input [3:0] S;
	output reg [15:0] O;
	
	always @(S)
	begin
		O = 16'b0;
		case({S})
			4'b0000: O[0]=1'b1;
			4'b0001: O[1]=1'b1;
			4'b0010: O[2]=1'b1;
			4'b0011: O[3]=1'b1;
			4'b0100: O[4]=1'b1;
			4'b0101: O[5]=1'b1;
			4'b0110: O[6]=1'b1;
			4'b0111: O[7]=1'b1;
			4'b1000: O[8]=1'b1;
			4'b1001: O[9]=1'b1;
			4'b1010: O[10]=1'b1;
			4'b1011: O[11]=1'b1;
			4'b1100: O[12]=1'b1;
			4'b1101: O[13]=1'b1;
			4'b1110: O[14]=1'b1;
			4'b1111: O[15]=1'b1;
		endcase
	end
endmodule