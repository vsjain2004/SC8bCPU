// Copyright (C) 2025  Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Altera and sold by Altera or its authorized distributors.  Please
// refer to the Altera Software License Subscription Agreements 
// on the Quartus Prime software download page.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 24.1std.0 Build 1077 03/04/2025 SC Lite Edition"
// CREATED		"Mon Oct  6 11:08:14 2025"

module CLA_8_bit(
	Cin,
	X,
	Y,
	Cout,
	Ov,
	S
);


input wire	Cin;
input wire	[7:0] X;
input wire	[7:0] Y;
output wire	Cout;
output wire	Ov;
output wire	[7:0] S;

wire	[7:0] S_ALTERA_SYNTHESIZED;
wire	[7:0] Z;
wire	SYNTHESIZED_WIRE_204;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_205;
wire	SYNTHESIZED_WIRE_206;
wire	SYNTHESIZED_WIRE_207;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_208;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_209;
wire	SYNTHESIZED_WIRE_210;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_211;
wire	SYNTHESIZED_WIRE_212;
wire	SYNTHESIZED_WIRE_213;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_214;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_215;
wire	SYNTHESIZED_WIRE_216;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_98;
wire	SYNTHESIZED_WIRE_217;
wire	SYNTHESIZED_WIRE_218;
wire	SYNTHESIZED_WIRE_136;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_138;
wire	SYNTHESIZED_WIRE_139;
wire	SYNTHESIZED_WIRE_140;
wire	SYNTHESIZED_WIRE_141;
wire	SYNTHESIZED_WIRE_142;
wire	SYNTHESIZED_WIRE_219;
wire	SYNTHESIZED_WIRE_188;
wire	SYNTHESIZED_WIRE_189;
wire	SYNTHESIZED_WIRE_190;
wire	SYNTHESIZED_WIRE_191;
wire	SYNTHESIZED_WIRE_192;
wire	SYNTHESIZED_WIRE_193;
wire	SYNTHESIZED_WIRE_194;
wire	SYNTHESIZED_WIRE_195;
wire	[7:0] SYNTHESIZED_WIRE_196;
wire	SYNTHESIZED_WIRE_197;
wire	SYNTHESIZED_WIRE_198;
wire	SYNTHESIZED_WIRE_199;
wire	SYNTHESIZED_WIRE_200;
wire	SYNTHESIZED_WIRE_202;

assign	Cout = SYNTHESIZED_WIRE_200;



assign	SYNTHESIZED_WIRE_206 = X[0] & Z[0];

assign	SYNTHESIZED_WIRE_202 = Cin & SYNTHESIZED_WIRE_204;

assign	SYNTHESIZED_WIRE_205 = Z[1] | X[1];

assign	SYNTHESIZED_WIRE_208 = Z[2] | X[2];

assign	SYNTHESIZED_WIRE_213 = Z[3] | X[3];

assign	SYNTHESIZED_WIRE_211 = Z[4] | X[4];

assign	SYNTHESIZED_WIRE_217 = Z[6] | X[6];

assign	SYNTHESIZED_WIRE_215 = Z[5] | X[5];


XOR_3_bit	b2v_inst16(
	.In1(X[0]),
	.In2(Z[0]),
	.In3(Cin),
	.Out(S_ALTERA_SYNTHESIZED[0]));


XOR_3_bit	b2v_inst17(
	.In1(X[1]),
	.In2(Z[1]),
	.In3(SYNTHESIZED_WIRE_1),
	.Out(S_ALTERA_SYNTHESIZED[1]));


XOR_3_bit	b2v_inst18(
	.In1(X[2]),
	.In2(Z[2]),
	.In3(SYNTHESIZED_WIRE_2),
	.Out(S_ALTERA_SYNTHESIZED[2]));


XOR_3_bit	b2v_inst19(
	.In1(X[3]),
	.In2(Z[3]),
	.In3(SYNTHESIZED_WIRE_3),
	.Out(S_ALTERA_SYNTHESIZED[3]));

assign	SYNTHESIZED_WIRE_14 = SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_206;


XOR_3_bit	b2v_inst20(
	.In1(X[7]),
	.In2(Z[7]),
	.In3(SYNTHESIZED_WIRE_207),
	.Out(S_ALTERA_SYNTHESIZED[7]));


XOR_3_bit	b2v_inst21(
	.In1(X[5]),
	.In2(Z[5]),
	.In3(SYNTHESIZED_WIRE_7),
	.Out(S_ALTERA_SYNTHESIZED[5]));


XOR_3_bit	b2v_inst22(
	.In1(X[4]),
	.In2(Z[4]),
	.In3(SYNTHESIZED_WIRE_8),
	.Out(S_ALTERA_SYNTHESIZED[4]));

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_204 & Cin;

assign	SYNTHESIZED_WIRE_22 = SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_204 & Cin;

assign	SYNTHESIZED_WIRE_2 = SYNTHESIZED_WIRE_14 | SYNTHESIZED_WIRE_15 | SYNTHESIZED_WIRE_209;

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_206 & SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_208;

assign	SYNTHESIZED_WIRE_3 = SYNTHESIZED_WIRE_210 | SYNTHESIZED_WIRE_21 | SYNTHESIZED_WIRE_22 | SYNTHESIZED_WIRE_23;


XOR_3_bit	b2v_inst28(
	.In1(X[6]),
	.In2(Z[6]),
	.In3(SYNTHESIZED_WIRE_24),
	.Out(S_ALTERA_SYNTHESIZED[6]));

assign	SYNTHESIZED_WIRE_62 = SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_212;

assign	SYNTHESIZED_WIRE_209 = X[1] & Z[1];

assign	SYNTHESIZED_WIRE_48 = SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_206;

assign	SYNTHESIZED_WIRE_47 = SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_209;

assign	SYNTHESIZED_WIRE_63 = SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_209;

assign	SYNTHESIZED_WIRE_61 = SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_210;


AND_5_bit	b2v_inst34(
	.In1(SYNTHESIZED_WIRE_213),
	.In2(SYNTHESIZED_WIRE_208),
	.In3(SYNTHESIZED_WIRE_205),
	.In4(SYNTHESIZED_WIRE_204),
	.In5(Cin),
	.Out(SYNTHESIZED_WIRE_49));


OR_5_bit	b2v_inst35(
	.In1(SYNTHESIZED_WIRE_212),
	.In2(SYNTHESIZED_WIRE_46),
	.In3(SYNTHESIZED_WIRE_47),
	.In4(SYNTHESIZED_WIRE_48),
	.In5(SYNTHESIZED_WIRE_49),
	.Out(SYNTHESIZED_WIRE_8));

assign	SYNTHESIZED_WIRE_65 = SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_204 & Cin;


AND_5_bit	b2v_inst37(
	.In1(SYNTHESIZED_WIRE_211),
	.In2(SYNTHESIZED_WIRE_213),
	.In3(SYNTHESIZED_WIRE_208),
	.In4(SYNTHESIZED_WIRE_205),
	.In5(SYNTHESIZED_WIRE_206),
	.Out(SYNTHESIZED_WIRE_64));

assign	SYNTHESIZED_WIRE_214 = X[4] & Z[4];

assign	SYNTHESIZED_WIRE_7 = SYNTHESIZED_WIRE_214 | SYNTHESIZED_WIRE_61 | SYNTHESIZED_WIRE_62 | SYNTHESIZED_WIRE_63 | SYNTHESIZED_WIRE_64 | SYNTHESIZED_WIRE_65;

assign	SYNTHESIZED_WIRE_210 = X[2] & Z[2];


AND_7_bit	b2v_inst40(
	.In1(SYNTHESIZED_WIRE_215),
	.In2(SYNTHESIZED_WIRE_211),
	.In3(SYNTHESIZED_WIRE_213),
	.In4(SYNTHESIZED_WIRE_208),
	.In5(SYNTHESIZED_WIRE_205),
	.In6(SYNTHESIZED_WIRE_204),
	.In7(Cin),
	.Out(SYNTHESIZED_WIRE_98));

assign	SYNTHESIZED_WIRE_97 = SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_206;


AND_5_bit	b2v_inst42(
	.In1(SYNTHESIZED_WIRE_215),
	.In2(SYNTHESIZED_WIRE_211),
	.In3(SYNTHESIZED_WIRE_213),
	.In4(SYNTHESIZED_WIRE_208),
	.In5(SYNTHESIZED_WIRE_209),
	.Out(SYNTHESIZED_WIRE_96));

assign	SYNTHESIZED_WIRE_93 = SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_214;

assign	SYNTHESIZED_WIRE_95 = SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_210;

assign	SYNTHESIZED_WIRE_94 = SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_212;

assign	SYNTHESIZED_WIRE_216 = X[5] & Z[5];


OR_7_bit	b2v_inst47(
	.In1(SYNTHESIZED_WIRE_216),
	.In2(SYNTHESIZED_WIRE_93),
	.In3(SYNTHESIZED_WIRE_94),
	.In4(SYNTHESIZED_WIRE_95),
	.In5(SYNTHESIZED_WIRE_96),
	.In6(SYNTHESIZED_WIRE_97),
	.In7(SYNTHESIZED_WIRE_98),
	.Out(SYNTHESIZED_WIRE_24));

assign	SYNTHESIZED_WIRE_142 = SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_204 & SYNTHESIZED_WIRE_205 & Cin & SYNTHESIZED_WIRE_208;


AND_7_bit	b2v_inst49(
	.In1(SYNTHESIZED_WIRE_217),
	.In2(SYNTHESIZED_WIRE_215),
	.In3(SYNTHESIZED_WIRE_211),
	.In4(SYNTHESIZED_WIRE_213),
	.In5(SYNTHESIZED_WIRE_208),
	.In6(SYNTHESIZED_WIRE_205),
	.In7(SYNTHESIZED_WIRE_206),
	.Out(SYNTHESIZED_WIRE_141));

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_209 & SYNTHESIZED_WIRE_208;

assign	SYNTHESIZED_WIRE_139 = SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_209;


AND_5_bit	b2v_inst51(
	.In1(SYNTHESIZED_WIRE_217),
	.In2(SYNTHESIZED_WIRE_215),
	.In3(SYNTHESIZED_WIRE_211),
	.In4(SYNTHESIZED_WIRE_213),
	.In5(SYNTHESIZED_WIRE_210),
	.Out(SYNTHESIZED_WIRE_140));

assign	SYNTHESIZED_WIRE_137 = SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_216;

assign	SYNTHESIZED_WIRE_138 = SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_212;

assign	SYNTHESIZED_WIRE_136 = SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_214;

assign	SYNTHESIZED_WIRE_218 = X[6] & Z[6];

assign	SYNTHESIZED_WIRE_207 = SYNTHESIZED_WIRE_218 | SYNTHESIZED_WIRE_136 | SYNTHESIZED_WIRE_137 | SYNTHESIZED_WIRE_138 | SYNTHESIZED_WIRE_139 | SYNTHESIZED_WIRE_140 | SYNTHESIZED_WIRE_141 | SYNTHESIZED_WIRE_142;

assign	SYNTHESIZED_WIRE_197 = SYNTHESIZED_WIRE_219 & SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_204 & SYNTHESIZED_WIRE_213;

assign	SYNTHESIZED_WIRE_195 = SYNTHESIZED_WIRE_219 & SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_205 & SYNTHESIZED_WIRE_208 & SYNTHESIZED_WIRE_206 & SYNTHESIZED_WIRE_213;


AND_7_bit	b2v_inst59(
	.In1(SYNTHESIZED_WIRE_219),
	.In2(SYNTHESIZED_WIRE_217),
	.In3(SYNTHESIZED_WIRE_215),
	.In4(SYNTHESIZED_WIRE_211),
	.In5(SYNTHESIZED_WIRE_213),
	.In6(SYNTHESIZED_WIRE_208),
	.In7(SYNTHESIZED_WIRE_209),
	.Out(SYNTHESIZED_WIRE_194));

assign	SYNTHESIZED_WIRE_46 = SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_210;

assign	SYNTHESIZED_WIRE_192 = SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_219 & SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_211 & SYNTHESIZED_WIRE_213 & SYNTHESIZED_WIRE_210;


AND_5_bit	b2v_inst61(
	.In1(SYNTHESIZED_WIRE_219),
	.In2(SYNTHESIZED_WIRE_217),
	.In3(SYNTHESIZED_WIRE_215),
	.In4(SYNTHESIZED_WIRE_211),
	.In5(SYNTHESIZED_WIRE_212),
	.Out(SYNTHESIZED_WIRE_193));

assign	SYNTHESIZED_WIRE_190 = SYNTHESIZED_WIRE_219 & SYNTHESIZED_WIRE_218;

assign	SYNTHESIZED_WIRE_191 = SYNTHESIZED_WIRE_219 & SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_215 & SYNTHESIZED_WIRE_214;

assign	SYNTHESIZED_WIRE_189 = SYNTHESIZED_WIRE_219 & SYNTHESIZED_WIRE_217 & SYNTHESIZED_WIRE_216;

assign	SYNTHESIZED_WIRE_219 = Z[7] | X[7];

assign	SYNTHESIZED_WIRE_188 = X[7] & Z[7];

assign	SYNTHESIZED_WIRE_198 = SYNTHESIZED_WIRE_188 | SYNTHESIZED_WIRE_189 | SYNTHESIZED_WIRE_190 | SYNTHESIZED_WIRE_191 | SYNTHESIZED_WIRE_192 | SYNTHESIZED_WIRE_193 | SYNTHESIZED_WIRE_194 | SYNTHESIZED_WIRE_195;


bit_1_to_8	b2v_inst68(
	.In(Cin),
	.Out(SYNTHESIZED_WIRE_196));


XOR_8_bit	b2v_inst69(
	.Control(SYNTHESIZED_WIRE_196),
	.In(Y),
	.Out(Z));

assign	SYNTHESIZED_WIRE_212 = X[3] & Z[3];

assign	SYNTHESIZED_WIRE_199 = SYNTHESIZED_WIRE_197 & Cin;

assign	SYNTHESIZED_WIRE_200 = SYNTHESIZED_WIRE_198 | SYNTHESIZED_WIRE_199;

assign	Ov = SYNTHESIZED_WIRE_200 ^ SYNTHESIZED_WIRE_207;

assign	SYNTHESIZED_WIRE_204 = Z[0] | X[0];

assign	SYNTHESIZED_WIRE_1 = SYNTHESIZED_WIRE_202 | SYNTHESIZED_WIRE_206;

assign	S = S_ALTERA_SYNTHESIZED;

endmodule
