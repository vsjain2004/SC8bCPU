module Control(
 input NOOP, IN, OUT, I_END, LDM, LDD, LDI, LDX, SWAP, STO, STI, STX, ADDM, ADDD, ADDI, ADDX, SUBM, SUBD, SUBI, SUBX, INC, DEC, LSL, LSR, ADDR, SUBR, MOV, CMP, CMD, CMI, CMX, SWAPR, JMP, JPN, JPE, JGT, JGE, ANDM, ANDD, ANDI, ANDX, ORM, ORD, ORI, ORX, XORM, XORD, XORI, XORX, NOT, ASR, CSL, CSR,
 input [1:0] RX, RY,
 input NF, OF, ZF,
 output REG_WLINE_1, REG_WLINE_0, REG_W_EN, REG_W_ADD_1, REG_W_ADD_0, REG_ADD_4, REG_ADD_3, REG_ADD_2, REG_ADD_1, REG_ADD_0, ADD_SUB, ALU_S_0, ALU_S_1, FLAG_W, ALU_SL_1, ALU_SL_0, DMEM_W_EN, DMEM_S_ADD, PC_LD_EN, PC_EN, OUT_EN, X_SEL, I_SEL, SWAP_R, ALU_S_2
 );

wire SYNTHESIZED_WIRE_0;
wire SYNTHESIZED_WIRE_1;
wire SYNTHESIZED_WIRE_2;
wire SYNTHESIZED_WIRE_3;
wire SYNTHESIZED_WIRE_5;
wire SYNTHESIZED_WIRE_6;
wire SYNTHESIZED_WIRE_8;
wire SYNTHESIZED_WIRE_9;
wire SYNTHESIZED_WIRE_10;
wire SYNTHESIZED_WIRE_11;
wire SYNTHESIZED_WIRE_12;
wire SYNTHESIZED_WIRE_13;
wire SYNTHESIZED_WIRE_14;
wire SYNTHESIZED_WIRE_15;
wire SYNTHESIZED_WIRE_20;
wire SYNTHESIZED_WIRE_21;
wire SYNTHESIZED_WIRE_22;
wire SYNTHESIZED_WIRE_23;
wire SYNTHESIZED_WIRE_24;
wire SYNTHESIZED_WIRE_25;
wire SYNTHESIZED_WIRE_26;
wire SYNTHESIZED_WIRE_27;
wire SYNTHESIZED_WIRE_28;
wire SYNTHESIZED_WIRE_29;
wire SYNTHESIZED_WIRE_30;
wire SYNTHESIZED_WIRE_31;
wire SYNTHESIZED_WIRE_34;
wire SYNTHESIZED_WIRE_35;
wire SYNTHESIZED_WIRE_36;
wire SYNTHESIZED_WIRE_37;

assign SYNTHESIZED_WIRE_0 = ADDI | CMI | SUBI | ANDI | ORI | XORI | LSL | LSR;

assign SYNTHESIZED_WIRE_1 = CMD | ANDM | CMX | ANDD | ORM | ANDX | ORD | ORX;

assign SYNTHESIZED_WIRE_2 = XORD | XORX | XORM | OUT | DEC | ASR | CSL | CSR;

assign SYNTHESIZED_WIRE_3 = ADDM | ADDX | ADDD | SUBM | SUBX | SUBD | INC | CMP;

assign SYNTHESIZED_WIRE_5 = SYNTHESIZED_WIRE_34 & RX[1];

assign SYNTHESIZED_WIRE_6 = MOV & RY[1];

assign SYNTHESIZED_WIRE_8 = SYNTHESIZED_WIRE_34 & RX[0];

assign SYNTHESIZED_WIRE_9 = MOV & RY[0];

assign SYNTHESIZED_WIRE_10 = SUBM | SUBX | SUBD | INC | CMP | CMD;

assign SYNTHESIZED_WIRE_11 = SUBI | CMI | ADDI | CMX | ADDR | SUBR;

assign SYNTHESIZED_WIRE_12 = ADDM | ADDX | ADDD | SUBM | SUBX | SUBD | CMP | CMD;

assign SYNTHESIZED_WIRE_13 = ANDM | ORM | ANDD | ORD | XORM | XORD | LSL | LSR;

assign SYNTHESIZED_WIRE_14 = ADDI | CMI | SUBI | ANDI | ORI | XORI | CSL | CSR;

assign SYNTHESIZED_WIRE_15 = LDX | ADDM | STX | ADDD | SUBD | SUBM | CMP | CMD;

assign SYNTHESIZED_WIRE_20 = SYNTHESIZED_WIRE_35 & JPN;

assign SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_36 & JGE;

assign SYNTHESIZED_WIRE_22 = SYNTHESIZED_WIRE_35 & SYNTHESIZED_WIRE_36 & JGT;

assign SYNTHESIZED_WIRE_23 = LDI | SUBI | ADDI | ANDI | ORI | XORI | SWAP | NOT;

assign SYNTHESIZED_WIRE_24 = SYNTHESIZED_WIRE_29 | SYNTHESIZED_WIRE_30 | XORX | SYNTHESIZED_WIRE_31;

assign SYNTHESIZED_WIRE_25 = SYNTHESIZED_WIRE_20 | SYNTHESIZED_WIRE_21 | JMP | SYNTHESIZED_WIRE_22;

assign SYNTHESIZED_WIRE_26 = ZF & JPE;

assign SYNTHESIZED_WIRE_27 = ADDI | CMI | SUBI | ANDI | ORI | XORI;

assign SYNTHESIZED_WIRE_28 = ADDD | INC | SUBD | MOV | ANDD | CMD | ORD | XORD;

assign SYNTHESIZED_WIRE_29 = LDM | LDX | LDD | ADDM | ADDX | ADDD | SUBM | SUBD;

assign SYNTHESIZED_WIRE_30 = ORD | XORM | XORD | ORX;

assign SYNTHESIZED_WIRE_31 = SUBX | MOV | INC | IN | ANDD | ANDM | ANDX | ORM;

assign SYNTHESIZED_WIRE_34 = SYNTHESIZED_WIRE_0 | SYNTHESIZED_WIRE_1 | SYNTHESIZED_WIRE_2 | SYNTHESIZED_WIRE_3 | ADDR | SUBR | SWAPR | NOT;

assign SYNTHESIZED_WIRE_35 =  ~ZF;

assign SYNTHESIZED_WIRE_36 = NF ~^ OF;

assign SYNTHESIZED_WIRE_37 = STI | STX | STO | SWAP;

assign REG_WLINE_1 = LDD | LDX | IN | LDI | SWAP;

assign REG_WLINE_0 = IN | LDM;

assign REG_W_EN = SYNTHESIZED_WIRE_23 | SYNTHESIZED_WIRE_24 | DEC | LSL | LSR | ASR | CSL | CSR;

assign REG_W_ADD_1 = RX[1];

assign REG_W_ADD_0 = RX[0];

assign REG_ADD_4 = INC | DEC;

assign REG_ADD_3 = (SYNTHESIZED_WIRE_37 & RX[1]) | ((ADDR | SUBR | SWAPR) & RY[1]);

assign REG_ADD_2 = (SYNTHESIZED_WIRE_37 & RX[0]) | ((ADDR | SUBR | SWAPR) & RY[0]);

assign REG_ADD_1 = SYNTHESIZED_WIRE_5 | LDX | STX | SYNTHESIZED_WIRE_6; //

assign REG_ADD_0 = SYNTHESIZED_WIRE_8 | LDX | STX | SYNTHESIZED_WIRE_9; //

assign ADD_SUB = SYNTHESIZED_WIRE_10 | SUBI | CMI | CMX | SUBR;

assign ALU_S_2 = LSL | LSR | NOT | ASR | CSL | CSR;

assign ALU_S_1 = ORM | ORI | ORD | ORX | XORD | XORM | XORI | XORX | ASR | CSL | CSR;

assign ALU_S_0 = ANDM | ANDI | ANDD | ANDX | XORD | XORM | XORI | XORX | LSL | LSR | CSL | CSR;

assign FLAG_W = SYNTHESIZED_WIRE_11 | SYNTHESIZED_WIRE_12;

assign ALU_SL_1 = SYNTHESIZED_WIRE_13 | SYNTHESIZED_WIRE_14 | SYNTHESIZED_WIRE_15 | ASR;

assign ALU_SL_0 = SYNTHESIZED_WIRE_27 | SYNTHESIZED_WIRE_28 | DEC;

assign DMEM_W_EN = STI | STX | STO | SWAP;

assign DMEM_S_ADD = STX | LDX;

assign PC_LD_EN = SYNTHESIZED_WIRE_25 | SYNTHESIZED_WIRE_26;

assign PC_EN =  ~I_END;

assign OUT_EN = OUT;

assign X_SEL = ADDX | CMX | SUBX | ANDX | ORX | XORX;

assign I_SEL = LDI | ADDI | STI | SUBI | ANDI | CMI | ORI | XORI;

assign SWAP_R = SWAPR;

endmodule
