module Zeros(Z);
	output [7:0] Z;

	assign Z = 8'b00000000;
endmodule