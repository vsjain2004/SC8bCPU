module Ones(O);
	output [7:0] O;

	assign O = 8'b11111111;
endmodule